library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package ethernet_rx_pkg is

end package ethernet_rx_pkg;

package body ethernet_rx_pkg is

end package body ethernet_rx_pkg;
